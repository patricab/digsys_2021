entity dff is
  port (
    clk     : in  std_logic;
    d       : in  std_logic;
    q       : out std_logic);
end dff;