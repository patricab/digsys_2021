-- p and q are large primes
-- n = p * q
-- C = M^e
-- M = C^d

M := 50

M^e mod n

C := 1
P := M

for i=0 to k-1
	if ei = 1
		C := C*P
	P := P*P
return C



A * B mod n

P = 0
for i=0 to k-1
	P = 2*P + A*B[k1-i]
	if P >= N
		P = P - N
	if P >= N
		P = P - N
	return P