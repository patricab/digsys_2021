entity mux2x1 is
  port (
    a       : in  std_logic;
    b       : in  std_logic;
    sel     : in  std_logic;
    y       : out std_logic);
end mux2x1;