package RSA is
   type states is (RSET, IDLE, PREP, CALC, FLIP, FNSH);
end package;

-- package body mary is
-- end package body;
